`timescale 1ns / 1ps
module uar_fsm_tb;
    logic clk;
    logic rst;
    logic sig;
    logic [161:0] data;
    logic ready;

    uar_fsm uar    (    .clk_in(clk),
                        .rst_in(rst),
                        .sig_in(sig),
                        .data_out(data),
                        .ready(ready));
    always begin
        #5;
        clk = !clk;
     end

     initial begin
        clk = 0;
        rst = 0;
        sig = 1;
        #10000;
        rst = 1;
        #10;
        rst = 0;
        
        #10;
        sig = 0;
        #104167;
        sig = 1;
        #104167;
        sig = 0;
        #104167;
        sig = 1;
        #104167;
        sig = 0;
        #104167;
        sig = 0;
        #104167;
        sig = 0;
        #104167;
        sig = 1;
        #104167;
        sig = 1;
        #104167;
        sig = 1;
        #104167;
        sig = 0;
        #104167;
        sig = 1;
        
        #2500000;
        
        sig = 0;
        #104167;
        sig = 1;
        #104167;
        sig = 0;
        #104167;
        sig = 1;
        #104167;
        sig = 0;
        #104167;
        sig = 0;
        #104167;
        sig = 0;
        #104167;
        sig = 1;
        #104167;
        sig = 1;
        #104167;
        sig = 1;
        #104167;
        sig = 0;
        #104167;
        sig = 1;
        #30000000;
        
        //Actual Transmission
        #10;
        sig = 0;
        #104167;
        sig = 1;
        #104167;
        sig = 0;
        #104167;
        sig = 1;
        #104167;
        sig = 0;
        #104167;
        sig = 1;
        #104167;
        sig = 0;
        #104167;
        sig = 1;
        #104167;
        sig = 0;
        #104167;
        sig = 1;
        #104167;
        sig = 0;
        #104167;
        sig = 1;
        #104167;
        sig = 0;
        #104167;
        sig = 1;
        #104167;
        sig = 0;
        #104167;
        sig = 1;
        #104167;
        sig = 0;
        #104167;
        sig = 1;
        #104167;
        
        sig = 0;
        #104167;
        sig = 1;
        #104167;
        sig = 0;
        #104167;
        sig = 1;
        #104167;
        sig = 0;
        #104167;
        sig = 1;
        #104167;
        sig = 0;
        #104167;
        sig = 1;
        #104167;
        sig = 0;
        #104167;
        sig = 1;
        #104167;
        sig = 0;
        #104167;
        sig = 1;
        #104167;
        sig = 0;
        #104167;
        sig = 1;
        #104167;
        sig = 0;
        #104167;
        sig = 1;
        #104167;
        sig = 0;
        #104167;
        sig = 1;
        #104167;
        
        sig = 0;
        #104167;
        sig = 1;
        #104167;
        sig = 0;
        #104167;
        sig = 1;
        #104167;
        sig = 0;
        #104167;
        sig = 1;
        #104167;
        sig = 0;
        #104167;
        sig = 1;
        #104167;
        sig = 0;
        #104167;
        sig = 1;
        #104167;
        sig = 0;
        #104167;
        sig = 1;
        #104167;
        sig = 0;
        #104167;
        sig = 1;
        #104167;
        sig = 0;
        #104167;
        sig = 1;
        #104167;
        sig = 0;
        #104167;
        sig = 1;
        #104167;
        
        sig = 0;
        #104167;
        sig = 1;
        #104167;
        sig = 0;
        #104167;
        sig = 1;
        #104167;
        sig = 0;
        #104167;
        sig = 1;
        #104167;
        sig = 0;
        #104167;
        sig = 1;
        #104167;
        sig = 0;
        #104167;
        sig = 1;
        #104167;
        sig = 0;
        #104167;
        sig = 1;
        #104167;
        sig = 0;
        #104167;
        sig = 1;
        #104167;
        sig = 0;
        #104167;
        sig = 1;
        #104167;
        sig = 0;
        #104167;
        sig = 1;
        #104167;
        
        sig = 0;
        #104167;
        sig = 1;
        #104167;
        sig = 0;
        #104167;
        sig = 1;
        #104167;
        sig = 0;
        #104167;
        sig = 1;
        #104167;
        sig = 0;
        #104167;
        sig = 1;
        #104167;
        sig = 0;
        #104167;
        sig = 1;
        #104167;
        sig = 0;
        #104167;
        sig = 1;
        #104167;
        sig = 0;
        #104167;
        sig = 1;
        #104167;
        sig = 0;
        #104167;
        sig = 1;
        #104167;
        sig = 0;
        #104167;
        sig = 1;
        #104167;
        
        sig = 0;
        #104167;
        sig = 1;
        #104167;
        sig = 0;
        #104167;
        sig = 1;
        #104167;
        sig = 0;
        #104167;
        sig = 1;
        #104167;
        sig = 0;
        #104167;
        sig = 1;
        #104167;
        sig = 0;
        #104167;
        sig = 1;
        #104167;
        sig = 0;
        #104167;
        sig = 1;
        #104167;
        sig = 0;
        #104167;
        sig = 1;
        #104167;
        sig = 0;
        #104167;
        sig = 1;
        #104167;
        sig = 0;
        #104167;
        sig = 1;
        #104167;
        
        sig = 0;
        #104167;
        sig = 1;
        #104167;
        sig = 0;
        #104167;
        sig = 1;
        #104167;
        sig = 0;
        #104167;
        sig = 1;
        #104167;
        sig = 0;
        #104167;
        sig = 1;
        #104167;
        sig = 0;
        #104167;
        sig = 1;
        #104167;
        sig = 0;
        #104167;
        sig = 1;
        #104167;
        sig = 0;
        #104167;
        sig = 1;
        #104167;
        sig = 0;
        #104167;
        sig = 1;
        #104167;
        sig = 0;
        #104167;
        sig = 1;
        #104167;
        
        sig = 0;
        #104167;
        sig = 1;
        #104167;
        sig = 0;
        #104167;
        sig = 1;
        #104167;
        sig = 0;
        #104167;
        sig = 1;
        #104167;
        sig = 0;
        #104167;
        sig = 1;
        #104167;
        sig = 0;
        #104167;
        sig = 1;
        #104167;
        sig = 0;
        #104167;
        sig = 1;
        #104167;
        sig = 0;
        #104167;
        sig = 1;
        #104167;
        sig = 0;
        #104167;
        sig = 1;
        #104167;
        sig = 0;
        #104167;
        sig = 1;
        #104167;
        
        sig = 0;
        #104167;
        sig = 1;
        #104167;
        sig = 0;
        #104167;
        sig = 1;
        #104167;
        sig = 0;
        #104167;
        sig = 1;
        #104167;
        sig = 0;
        #104167;
        sig = 1;
        #104167;
        sig = 0;
        #104167;
        sig = 1;
        #104167;
        sig = 0;
        #104167;
        sig = 1;
        #104167;
        sig = 0;
        #104167;
        sig = 1;
        #104167;
        sig = 0;
        #104167;
        sig = 1;
        #104167;
        sig = 0;
        #104167;
        sig = 1;
        //Whole Board
        
        #10000000;
        
     end
endmodule
